module ID_EX(Clk,Reset,Flush,ControlsIn,Data1_In,Data2_In,JEQAddrIn,JMPAddrIn,Imm8In,Reg1In,Reg2In,
