module IMEM(Addr,Ins);
input[15:0]Addr;
output[15:0]Ins;

wire[15:0]ROM[29:0];
assign Ins=ROM[Addr];
assign ROM[0]=16'b0001100000001010;//MOVI,R0,10
assign ROM[1]=16'b0000000000000000;
assign ROM[2]=16'b0000000000000000;
assign ROM[3]=16'b0001100100001110;//MOVI,R0,14
assign ROM[4]=16'b0000100000100000;//ADD,R0,R1
assign ROM[5]=16'b0000000000000000;
assign ROM[6]=16'b0000000000000000;
assign ROM[7]=16'b0001101000000100;//MOVI,R2,4
assign ROM[8]=16'b0001000001000000;//SUB,R0,R2
assign ROM[9]=16'b0000000000000000;//NOP
assign ROM[10]=16'b0000000000000000;//NOP
assign ROM[11]=16'b0001101100000000;//MOVI,R3,0
assign ROM[12]=16'b0000000000000000;//NOP
assign ROM[13]=16'b0000000000000000;//NOP
assign ROM[14]=16'b0000000000000000;//NOP
assign ROM[15]=16'b0010100001100000;//STO,R0,R3 MEM[0]=20
assign ROM[16]=16'b0000101101000000;//ADD,R3,R2 R3=4
assign ROM[17]=16'b0001110000010000;//MOVI,R4,16
assign ROM[18]=16'b0000000000000000;//NOP
assign ROM[19]=16'b0000000000000000;//NOP
assign ROM[20]=16'b0000000000000000;//NOP
assign ROM[21]=16'b0011100010001000;//JEQ,R0,R4,8
assign ROM[22]=16'b0000110001000000;//ADD,R4,R2
assign ROM[23]=16'b0001110100000000;//MOVI,R5,0
assign ROM[24]=16'b0000000000000000;//NOP
assign ROM[25]=16'b0000000000000000;//NOP
assign ROM[26]=16'b0000000000000000;//NOP
assign ROM[27]=16'b0010011010100000;//LODR R6,R5 R6=Mem[0]=20
assign ROM[28]=16'b0011011111111001;//JMP -7
assign ROM[29]=16'b0000110101000000;//ADD,R5,R2
endmodule
